module multiplier_tb_2();

reg [31: 0]in_data_A;
reg [31: 0]in_data_B;
wire[31: 0]out_data;

wire done = 0;
wire overflow_flag = 0;
wire underflow_flag = 0;



integer i;
integer failed_test_count;


localparam T = 150;

reg [511: 0] Data_to_input_A;
reg [511: 0] Data_to_input_B;
reg [511: 0] Expected_data;
reg [511: 0] Data_output;

multiplier #(32) inst (in_data_A,in_data_B,out_data,done, overflow_flag, underflow_flag);

initial begin
	Data_to_input_A <= 512'b00000000100000000000000000000000100000001000000000000000000000000111111101000000000010001000000001111111010000000000100010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000100000010100000000000000000000011000000101000000000000000000000001111110000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000100000011110100000000000000000001000001110010000000000000000000;
	Data_to_input_B <= 512'b00000001100000000000000000000000000000011000000000000000000000000111111101000011000010001000000011111111010000110000100010000000000000000000000000000000000000001000000000000000000000000000000001111111100000000000000000000000111111111000000000000000000000000100000011000000000000000000000001000000110000000000000000000000010000001100100000000000000000000111111110000000000000000000000010000000000000000000000000000000010000001111010000000000000000000000000000000000000000000000000001000000101000000000000000000000;
	Expected_data   <= 512'b0000000000000000000000000000000010000000000000000000000000000000011111111XXXXXXXXXXXXXXXXXXXXXXX111111111XXXXXXXXXXXXXXXXXXXXXXX00000000000000000000000000000000100000000000000000000000000000000111111110000000000000000000000011111111100000000000000000000000010000011111000000000000000000001100000111110000000000000000000001000000010010000000000000000000X11111111XXXXXXXXXXXXXXXXXXXXXXXX11111111XXXXXXXXXXXXXXXXXXXXXXX011111111000000000000000000000000000000000000000000000000000000001000010111110100000000000000000;
	
	for(i = 0; i< 512; i = i+32)
	begin
		#(T)
		$monitor ("%b      %b		%b\t",in_data_A,in_data_B,out_data);
		in_data_A = Data_to_input_A[i+:32];
		in_data_B = Data_to_input_B[i+:32];
		#(T)
		Data_output[i+:32] = out_data;
	end
	
		$display("output = %b", Data_output);
		failed_test_count =0;
		for(i = 0; i< 512; i = i+32)
		begin
			if(Data_output[i+:32] != Expected_data[i+:32]) begin
				$display("Test Input A: %b Test Input B: %b Expected Output: %b Actual Output: %b \n",Data_to_input_A[i+:32],Data_to_input_B[i+:32],Expected_data[i+:32],Data_output[i+:32]);
				failed_test_count = failed_test_count+1;
			end
		end
		if (failed_test_count ==0) $display("All Tests succeeded\n", i);
		else begin
			$display("failed test count: %d\n",failed_test_count);
		end
		
	$finish;
end
endmodule