module goldschmidtVersion2 (a,b,start,clk,clrn,q,busy,ready,yn);
input [31:0] a; // dividend: .1xxx...x
input [31:0] b; // divisor: .1xxx...x
input start; // start
input clk, clrn; // clock and reset
output [31:0] q; // quotient: x.xxx...x
output reg busy; // busy
output reg ready; // ready
//output [2:0] count; // counter
output [31:0] yn; // .11111...1
reg [63:0] reg_a; // x.xxxx...x
reg [63:0] reg_b; // 0.xxxx...x
reg [63:0] reg_b_Negative; // 0.xxxx...x
reg [2:0] count;
wire [63:0] two_minus_yi;// 2's complement
wire done,overflow,underflow;
wire mostSignificant1 = 32'b100000000000_0000000000000000000000000000000000000000000000000000;
wire [31:0] dNegative = q | mostSignificant1;
wire [31:0] twoWire = 32'b0_10000000000_0000000000000000000000000000000000000000000000000000;
wire [127:0] xi = reg_a * two_minus_yi; // 0x.xxx...x
wire [127:0] yi = reg_b * two_minus_yi; // 0x.xxx...x
//assign q = reg_a[63:32] + |reg_a[31:29]; // rounding up
assign q = reg_a[63:32];
assign yn = reg_b[62:31];
always @ (posedge clk or negedge clrn) begin
if (!clrn) begin
busy <= 0;
ready <= 0;
end else begin
if (start) begin
reg_a <= {1'b0,a,31'b0}; // 0.1x...x0...0
reg_b <= {1'b0,b,31'b0}; // 0.1x...x0...0
reg_b_Negative <= {1'b1,b,31'b0};
busy <= 1;
ready <= 0;
count <= 0;
end else begin
reg_a <= xi[126:63]; // x.xxx...x
reg_b <= yi[126:63]; // 0.xxx...x
reg_b_Negative <= reg_b | mostSignificant1;
count <= count + 3'b1; // count++
if (count == 3'h7) begin // finish
busy <= 0;
ready <= 1; // q is ready
end
end
end
end

adder #(32) inst (twoWire,reg_b_Negative,two_minus_yi,done,overflow,underflow);
//multiplier #(32) inst2 (reg_a,);

endmodule